module FNTT (
    input [63:0] data_in,
    input [7:0] omega,
    input [7:0] mod,
    input [7:0] N
    output [63:0] data_out
);

endmodule