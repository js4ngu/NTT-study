library verilog;
use verilog.vl_types.all;
entity reverse_bits_tb is
end reverse_bits_tb;
