library verilog;
use verilog.vl_types.all;
entity naiveNTT_tb is
end naiveNTT_tb;
