library verilog;
use verilog.vl_types.all;
entity bit_reverse_ordered_sv_unit is
end bit_reverse_ordered_sv_unit;
