library verilog;
use verilog.vl_types.all;
entity \_4point2dButterfly_sv_unit\ is
end \_4point2dButterfly_sv_unit\;
