library verilog;
use verilog.vl_types.all;
entity tb_fntt is
end tb_fntt;
