library verilog;
use verilog.vl_types.all;
entity \_16point2dButterfly_sv_unit\ is
end \_16point2dButterfly_sv_unit\;
