library verilog;
use verilog.vl_types.all;
entity tb_8point_BM is
end tb_8point_BM;
