module simpleNTT(a,o);
    input a[0:5][0:8];
    output o[0:5][0:8];

    
endmodule