library verilog;
use verilog.vl_types.all;
entity tb_4pont_BM is
end tb_4pont_BM;
