library verilog;
use verilog.vl_types.all;
entity dataslice_tb is
end dataslice_tb;
