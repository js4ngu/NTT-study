library verilog;
use verilog.vl_types.all;
entity tb_bit_reverse_ordered is
end tb_bit_reverse_ordered;
