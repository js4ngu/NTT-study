library verilog;
use verilog.vl_types.all;
entity omgea_genrator_sv_unit is
end omgea_genrator_sv_unit;
