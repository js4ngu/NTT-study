library verilog;
use verilog.vl_types.all;
entity tb_4vs8_CMP is
end tb_4vs8_CMP;
