library verilog;
use verilog.vl_types.all;
entity naiveNTTPolyMul_tb is
end naiveNTTPolyMul_tb;
