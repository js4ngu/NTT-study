library verilog;
use verilog.vl_types.all;
entity \_8point2dnaiveFNTT_sv_unit\ is
end \_8point2dnaiveFNTT_sv_unit\;
