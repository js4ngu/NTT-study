library verilog;
use verilog.vl_types.all;
entity naiveINTT_tb is
end naiveINTT_tb;
