`timescale 1ns/10ps

module naiveINTT_tb;
    reg [63:0] datain;
    wire [63:0] dataout;
    wire [63:0] result;
    reg [7:0] omega;
    reg [7:0] invOmega;
    reg [7:0] invN;
    reg [7:0] mod;

    initial begin
        mod = 17;
        omega = 9;
        invOmega = 2;
        invN = 15;
        //datain = 64'h03_01_02_06_00_00_00_00; //target
        datain = 64'h00_00_00_00_06_02_01_03; //target - Clear! ; output also reverse
        #10
        $finish;
    end
    naiveNTT u0 (
        .data_in(datain),
        .omega(omega),
        .mod(mod),
        .data_out(dataout)
    );

    naiveINTT u1(
        .data_in(dataout),
        .invN(invN),
        .invOmega(invOmega),
        .mod(mod),
        .data_out(result)
    );
endmodule


// 06  08 11 12  02  06 10  03

// 일단 in