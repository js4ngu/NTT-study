library verilog;
use verilog.vl_types.all;
entity tb_4piont_BM is
end tb_4piont_BM;
