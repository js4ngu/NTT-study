library verilog;
use verilog.vl_types.all;
entity tb_4point_BM is
end tb_4point_BM;
